module main;
initial
begin
    $display("Hello, World");
    #10 $finish;
end
endmodule
